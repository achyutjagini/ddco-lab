// Module 4-bit ripple carry adder


module fulladdR(input wire [3:0] a, b, input wire cin, output wire [3:0] sum, output wire cout);

  
 // Instantiate full adder modules here.

wire [2:0] c;
 
 fulladd u0 (                  );

  fulladd u1 (                 );

  fulladd u2 (                 );

  fulladd u3 (                 );


endmodule 


    

module mux4 (input wire [0:3] i, input wire j1, j0, output wire o);
 
 wire  t0, t1;
  
mux2 mux2_0 (                   );

  mux2 mux2_1 (                 );

  mux2 mux2_2 (                  );

endmodule


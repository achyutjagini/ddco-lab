module fulladd(input wire a, b, cin, output wire sum, cout);
wire [4:0] t;

   
 xor2 x0(               );

 xor2 x1(               );


 and2 a0(              );
  
 and2 a1(               );
   
 and2 a2(               );

    
  or2 o0(                    );
 
   or2 o1(                 );

endmodule
